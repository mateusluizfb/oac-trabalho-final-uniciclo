library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity mem_dados_tb is
end entity ; -- mem_dados_tb
architecture arch of mem_dados_tb is

begin

end architecture ; -- arch